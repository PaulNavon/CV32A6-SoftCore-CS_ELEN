/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_32 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 877;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00206567_616d6920,
        64'h746f6f62_20676e69,
        64'h79706f63_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_09202020,
        64'h20203a64_69756720,
        64'h6e6f6974_69747261,
        64'h70090a0d_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_093a6162,
        64'h6c20746e_65727275,
        64'h63090a0d_00000009,
        64'h3a646576_72657365,
        64'h72090a0d_00093a72,
        64'h65646165_685f6372,
        64'h63090a0d_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h003a7265_64616568,
        64'h20656c62_6174206e,
        64'h6f697469_74726170,
        64'h20747067_0000203a,
        64'h65756c61_76206e72,
        64'h75746572_2079706f,
        64'h63206473_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h0000000a_0d216465,
        64'h7a696c61_6974696e,
        64'h69206473_00000000,
        64'h0a0d676e_69746978,
        64'h65202e2e_2e647320,
        64'h657a696c_61697469,
        64'h6e692074_6f6e2064,
        64'h6c756f63_0000002e,
        64'h0000000a_0d6b636f,
        64'h6c622044_53206461,
        64'h65722074_6f6e2064,
        64'h6c756f63_0000000a,
        64'h0d202e2e_2e445320,
        64'h676e697a_696c6169,
        64'h74696e69_00000031,
        64'h34646d63_00000035,
        64'h35646d63_00000000,
        64'h30646d63_00000020,
        64'h3a206573_6e6f7073,
        64'h65720920_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000a0d_2164657a,
        64'h696c6169_74696e69,
        64'h20495053_00000a0d,
        64'h00007830_203a7375,
        64'h74617473_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_42424242,
        64'h0000000a_0000006f,
        64'h0000006c_00000061,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_68746469,
        64'h772d6f69_2d676572,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00736567_6e617200,
        64'h656c646e_61687000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_00687461,
        64'h702d7475_6f647473,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_006c6f72,
        64'h746e6f63_d8000000,
        64'h08000000_03000000,
        64'h02000000_0e010000,
        64'h04000000_03000000,
        64'h00100000_00000018,
        64'h67000000_08000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_1f010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h34010000_04000000,
        64'h03000000_02000000,
        64'h2a010000_04000000,
        64'h03000000_01000000,
        64'h1f010000_04000000,
        64'h03000000_02000000,
        64'h0e010000_04000000,
        64'h03000000_00c20100,
        64'h00010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000010_67000000,
        64'h08000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_f5000000,
        64'h04000000_03000000,
        64'h07000000_e2000000,
        64'h04000000_03000000,
        64'h00000004_0000000c,
        64'h67000000_08000000,
        64'h03000000_09000000,
        64'h01000000_0b000000,
        64'h01000000_c4000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_d8000000,
        64'h08000000_03000000,
        64'h00000c00_00000002,
        64'h67000000_08000000,
        64'h03000000_07000000,
        64'h01000000_03000000,
        64'h01000000_c4000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hbd000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h01000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_00000008,
        64'h00000080_67000000,
        64'h08000000_03000000,
        64'h00007972_6f6d656d,
        64'h5b000000_07000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6f6d656d_01000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'hb5000000_04000000,
        64'h03000000_00006374,
        64'h6e692d75_70632c76,
        64'h63736972_1b000000,
        64'h0f000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h85000000_00000000,
        64'h03000000_00003233,
        64'h76732c76_63736972,
        64'h7c000000_0b000000,
        64'h03000000_00616d69,
        64'h32337672_72000000,
        64'h08000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h01000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0c050000_41010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h44050000_38000000,
        64'h85060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0000006f_8dcff0ef,
        64'h80050513_00001517,
        64'h8e8ff0ef_80850513,
        64'h00001517_8f4ff0ef,
        64'h81050513_00001517,
        64'h900ff0ef_81850513,
        64'h00001517_90cff0ef,
        64'h82050513_00001517,
        64'h918ff0ef_81c50513,
        64'h00001517_8dcff0ef,
        64'h00112623_a0050513,
        64'h20058593_ff010113,
        64'h02626537_0001c5b7,
        64'hf11ff06f_ffe00493,
        64'h948ff0ef_88c50513,
        64'h00001517_a1cff0ef,
        64'h41f4d593_00048513,
        64'h960ff0ef_99050513,
        64'h00001517_96cff0ef,
        64'h98850513_00001517,
        64'hf49ff06f_ffe00493,
        64'h980ff0ef_8c450513,
        64'h00001517_a54ff0ef,
        64'h41fad593_000a8513,
        64'h998ff0ef_9c850513,
        64'h00001517_9a4ff0ef,
        64'h9c050513_00001517,
        64'hf81ff06f_ffe00493,
        64'h9b8ff0ef_8fc50513,
        64'h00001517_a8cff0ef,
        64'h41f4d593_00048513,
        64'h9d0ff0ef_a0050513,
        64'h00001517_9dcff0ef,
        64'h9f850513_00001517,
        64'hfb9ff06f_fff00493,
        64'h9f0ff0ef_9d050513,
        64'h00001517_00008067,
        64'h03010113_00812c03,
        64'h00c12b83_01012b03,
        64'h01412a83_01812a03,
        64'h01c12983_02012903,
        64'h02412483_02812403,
        64'h00048513_02c12083,
        64'hfd040113_a34ff0ef,
        64'hc0850513_00001517,
        64'h04051e63_00050493,
        64'hb91ff0ef_40b60633,
        64'h00160613_000b8513,
        64'h020c2583_028c2603,
        64'ha60ff0ef_c2050513,
        64'h00001517_f36a94e3,
        64'h080a0a13_08098993,
        64'h08048913_a7cff0ef,
        64'h001a8a93_9c450513,
        64'h00001517_ff249ae3,
        64'hbe4ff0ef_00148493,
        64'h0004c503_a9cff0ef,
        64'hc5050513_00001517,
        64'hb70ff0ef_0149a583,
        64'h0109a503_ab4ff0ef,
        64'hc5850513_00001517,
        64'hb88ff0ef_0089a503,
        64'h00c9a583_accff0ef,
        64'hc6050513_00001517,
        64'hba0ff0ef_fb890493,
        64'h0009a503_0049a583,
        64'hae8ff0ef_c6c50513,
        64'h00001517_ff349ae3,
        64'hc4cff0ef_00148493,
        64'h0004c503_000a0493,
        64'hb08ff0ef_c7050513,
        64'h00001517_ff449ae3,
        64'hc6cff0ef_00148493,
        64'h0004c503_f8090493,
        64'hb28ff0ef_c7450513,
        64'h00001517_c88ff0ef,
        64'h0ffaf513_b3cff0ef,
        64'hc7050513_00001517,
        64'h00400b13_01010a13,
        64'h02010993_08010913,
        64'h1a051663_00050a93,
        64'h00010c13_cadff0ef,
        64'h00100613_00010513,
        64'he0010113_04892583,
        64'hb78ff0ef_abc50513,
        64'h00001517_be4ff0ef,
        64'h05412503_b8cff0ef,
        64'hca050513_00001517,
        64'hbf8ff0ef_05012503,
        64'hba0ff0ef_c9450513,
        64'h00001517_c74ff0ef,
        64'h04812503_04c12583,
        64'hbb8ff0ef_c8c50513,
        64'h00001517_c8cff0ef,
        64'h02012503_02412583,
        64'hbd0ff0ef_c9450513,
        64'h00001517_ca4ff0ef,
        64'h01812503_01c12583,
        64'hbe8ff0ef_c9850513,
        64'h00001517_c54ff0ef,
        64'h01412503_bfcff0ef,
        64'hc9c50513_00001517,
        64'hc68ff0ef_01012503,
        64'hc10ff0ef_ca050513,
        64'h00001517_c7cff0ef,
        64'h00c12503_c24ff0ef,
        64'hca850513_00001517,
        64'hc90ff0ef_00812503,
        64'hc38ff0ef_cac50513,
        64'h00001517_d0cff0ef,
        64'h00012503_00412583,
        64'hc50ff0ef_cb450513,
        64'h00001517_c5cff0ef,
        64'hca450513_00001517,
        64'h2e051a63_00050493,
        64'h00010913_dbdff0ef,
        64'h00060593_00010513,
        64'he0010113_00100613,
        64'hc88ff0ef_c9050513,
        64'h00001517_28051e63,
        64'hc65ff0ef_00050b93,
        64'h03010413_01812423,
        64'h01612823_01512a23,
        64'h01412c23_01312e23,
        64'h03212023_02912223,
        64'h02112623_01712623,
        64'h02812423_fd010113,
        64'hfc1ff06f_fff00413,
        64'hcd8ff0ef_c9850513,
        64'h00001517_fe041ae3,
        64'hf6cff0ef_fff40413,
        64'h0ff00513_00800413,
        64'h00008067_0b010113,
        64'h09012b03_09c12983,
        64'h0a812403_00040513,
        64'h0ac12083_08812c03,
        64'h08c12b83_09412a83,
        64'h09812a03_0a012903,
        64'h0a412483_fb0ff0ef,
        64'h0ff00513_955ff0ef,
        64'h00c00513_00000593,
        64'h00100613_ffe00413,
        64'hfe5ff06f_d4cff0ef,
        64'hd2850513_00001517,
        64'h0180006f_00000413,
        64'hf1304ee3_fff98993,
        64'h00f98a63_035787b3,
        64'h40e787b3_4067d793,
        64'h41f9d713_034997b3,
        64'h02879e63_000c0b13,
        64'h0107d793_01079793,
        64'h012567b3_819ff0ef,
        64'h01095913_0ff00513,
        64'h01091913_00851913,
        64'h82dff0ef_0ff00513,
        64'hf92c14e3_04070b13,
        64'h040c0c13_fb6714e3,
        64'h01045413_00170713,
        64'h01041413_00f44433,
        64'h0177f7b3_00541793,
        64'h41045413_01041413,
        64'h00f44433_00c41793,
        64'h41045413_01041413,
        64'h00f44433_00f7f793,
        64'h00445793_00f44433,
        64'h0107d793_01079793,
        64'h00074403_0087e7b3,
        64'h00841413_00845793,
        64'h000c0713_959ff0ef,
        64'h00010513_04000593,
        64'h000c0613_00000413,
        64'h040b0b13_200c0913,
        64'h000b0c13_fe951ce3,
        64'h8c5ff0ef_0ff00513,
        64'h3e800a93_0fe00493,
        64'hdd3a0a13_fe0b8b93,
        64'h09812423_0b212023,
        64'h09512a23_0a912223,
        64'h00002bb7_10625a37,
        64'h09712623_09412c23,
        64'h18051263_a9dff0ef,
        64'h01200513_00100613,
        64'hfed79ae3_00478793,
        64'h08010693_00e7a023,
        64'hfff00713_00010793,
        64'h00060993_00050b13,
        64'h0a812423_0a112623,
        64'h09612823_09312e23,
        64'hf5010113_00008067,
        64'h01055513_01051513,
        64'h00f54533_00e7f7b3,
        64'h00551793_fe070713,
        64'h00002737_41055513,
        64'h01051513_00f54533,
        64'h00c51793_41055513,
        64'h01051513_00f5c533,
        64'h00f7f793_0045d793,
        64'h00f5c5b3_0107d793,
        64'h01079793_00a7e7b3,
        64'h00851513_00855793,
        64'h00008067_07f57513,
        64'h00f54533_0ff7f793,
        64'h00451793_00b54533,
        64'h00f54533_0045d513,
        64'h0075d793_00b575b3,
        64'hfc9ff06f_ffe00513,
        64'h00008067_01010113,
        64'hfff00513_00012903,
        64'h00412483_00812403,
        64'h00c12083_00008067,
        64'h01010113_00012903,
        64'h00412483_00812403,
        64'h00c12083_ffd57513,
        64'h40a00533_00153513,
        64'he7dff0ef_04050463,
        64'hd61ff0ef_f94ff0ef,
        64'hed850513_00001517,
        64'h8f5ff0ef_00090513,
        64'hfa8ff0ef_f2850513,
        64'h00001517_fb4ff0ef,
        64'hf4450513_00001517,
        64'hfc0ff0ef_f3450513,
        64'h00001517_fd241ee3,
        64'h06048863_a59ff0ef,
        64'h0ff00513_fff48493,
        64'h00050413_c05ff0ef,
        64'h00000513_00000593,
        64'h09500613_00100913,
        64'h71048493_000024b7,
        64'hfe041ae3_a89ff0ef,
        64'hfff40413_0ff00513,
        64'h00a00413_815ff0ef,
        64'hfbc50513_00001517,
        64'h9e1ff0ef_01212023,
        64'h00912223_00812423,
        64'h00112623_ff010113,
        64'h00008067_01010113,
        64'h00412483_00812403,
        64'h00143513_00c12083,
        64'hf4940ce3_ad9ff0ef,
        64'h0ff00513_85dff0ef,
        64'hfa050513_00001517,
        64'h9bdff0ef_00040513,
        64'h871ff0ef_ff050513,
        64'h00001517_87dff0ef,
        64'h01c50513_00001517,
        64'h889ff0ef_ffc50513,
        64'h00001517_00050413,
        64'hcb9ff0ef_02900513,
        64'h400005b7_07700613,
        64'h8a9ff0ef_fec50513,
        64'h00001517_a09ff0ef,
        64'h00040513_8bdff0ef,
        64'h03c50513_00001517,
        64'h8c9ff0ef_06050513,
        64'h00001517_8d5ff0ef,
        64'h04850513_00001517,
        64'hb65ff0ef_0ff00513,
        64'h00050413_d0dff0ef,
        64'h03700513_00000593,
        64'h06500613_00100493,
        64'h00812423_00112623,
        64'h00912223_ff010113,
        64'h00008067_01010113,
        64'h00153513_00812403,
        64'hfff40513_00c12083,
        64'h929ff0ef_06c50513,
        64'h00001517_a89ff0ef,
        64'h00040513_93dff0ef,
        64'h0bc50513_00001517,
        64'h949ff0ef_0e050513,
        64'h00001517_955ff0ef,
        64'h0c850513_00001517,
        64'hbe5ff0ef_0ff00513,
        64'h00050413_d8dff0ef,
        64'h00812423_00112623,
        64'h03700513_00000593,
        64'h06500613_ff010113,
        64'h00008067_01010113,
        64'h0017b513_00012903,
        64'h00412483_f5690793,
        64'h00812403_00c12083,
        64'hfe8792e3_00f4f793,
        64'h00008067_01010113,
        64'h00012903_00412483,
        64'h00812403_00c12083,
        64'h00f40e63_00000513,
        64'h00100793_c59ff0ef,
        64'h0ff00513_c61ff0ef,
        64'h0ff00513_00050913,
        64'hc6dff0ef_0ff00513,
        64'h00050493_c79ff0ef,
        64'h0ff00513_c81ff0ef,
        64'h0ff00513_c89ff0ef,
        64'h0ff00513_00050413,
        64'he31ff0ef_01212023,
        64'h00912223_00812423,
        64'h00112623_00800513,
        64'h1aa00593_08700613,
        64'hff010113_00008067,
        64'h01010113_00000513,
        64'h00012903_00412483,
        64'h00812403_00c12083,
        64'h00008067_01010113,
        64'h00012903_00090513,
        64'h00412483_00812403,
        64'h00c12083_a6dff0ef,
        64'h1b050513_00001517,
        64'hbcdff0ef_00090513,
        64'ha81ff0ef_20050513,
        64'h00001517_a8dff0ef,
        64'h21c50513_00001517,
        64'ha99ff0ef_20c50513,
        64'h00001517_fd241ee3,
        64'h04048e63_d31ff0ef,
        64'h0ff00513_fff48493,
        64'h00050413_eddff0ef,
        64'h00000513_00000593,
        64'h09500613_00100913,
        64'h71048493_00812423,
        64'h00112623_01212023,
        64'h000024b7_00912223,
        64'hff010113_aedff06f,
        64'h01010113_23450513,
        64'h00001517_00412483,
        64'h00c12083_00812403,
        64'hc5dff0ef_00040513,
        64'hb11ff0ef_29050513,
        64'h00001517_b1dff0ef,
        64'h00048513_b25ff0ef,
        64'h00058413_00812423,
        64'h00112623_2a450513,
        64'h00001517_00050493,
        64'h00912223_ff010113,
        64'h00008067_01010113,
        64'h00012903_00412483,
        64'h00812403_00c12083,
        64'hfe07c4e3_fff40413,
        64'h4187d793_01851793,
        64'hdf5ff0ef_0ff00513,
        64'h00040e63_0080006f,
        64'h06400413_e09ff0ef,
        64'h00048513_e11ff0ef,
        64'h0ff47513_e19ff0ef,
        64'h0ff57513_00845513,
        64'he25ff0ef_0ff57513,
        64'h01045513_e31ff0ef,
        64'h01845513_e39ff0ef,
        64'h04096513_e41ff0ef,
        64'h00060493_00058413,
        64'h00912223_00812423,
        64'h00112623_0ff00513,
        64'h00050913_01212023,
        64'hff010113_e69ff06f,
        64'h0ff00513_00008067,
        64'hfff00513_00008067,
        64'h00000513_06e7a023,
        64'h00600713_06d72823,
        64'h00070793_fff00693,
        64'h20000737_fec594e3,
        64'hfef60fa3_00160613,
        64'h0006a783_fe079ce3,
        64'h0017f793_00072783,
        64'h06c68693_06470713,
        64'h00b605b3_00070693,
        64'h20000737_00008067,
        64'h00000513_06e7a023,
        64'h00600713_06d72823,
        64'h00070793_fff00693,
        64'h20000737_02059263,
        64'hfe079ce3_0017f793,
        64'h00072783_06478713,
        64'h06d7a023_10600693,
        64'h200007b7_fe079ce3,
        64'hfff78793_00000013,
        64'h03200793_fed51ae3,
        64'h00f72023_00150513,
        64'h00054783_06870713,
        64'h00b506b3_20000737,
        64'h02058063_06e7a823,
        64'hffe00713_200007b7,
        64'h0cb7e863_10000793,
        64'hfadff06f_ccdff0ef,
        64'h41050513_00001517,
        64'hda1ff0ef_00000593,
        64'h00042503_ce5ff0ef,
        64'h44050513_00001517,
        64'h00008067_01010113,
        64'h00412483_0ff4f513,
        64'h06e7a023_00600713,
        64'h00070793_06d72823,
        64'hfff00693_00812403,
        64'h00c12083_20000737,
        64'h02078a63_0017f793,
        64'h00042783_06c7a483,
        64'h200007b7_fe079ce3,
        64'h0017f793_00042783,
        64'h06478413_06e7a023,
        64'h10600713_200007b7,
        64'hfe079ce3_fff78793,
        64'h00000013_06400793,
        64'h06a7a423_06d7a823,
        64'hffe00693_00912223,
        64'h00812423_00112623,
        64'h200007b7_ff010113,
        64'hd81ff06f_01010113,
        64'h4cc50513_00001517,
        64'h00012903_00412483,
        64'h00c12083_00812403,
        64'h06f42023_00600793,
        64'hda9ff0ef_4ec50513,
        64'h00001517_e7dff0ef,
        64'h00000593_00048513,
        64'hdc1ff0ef_4f850513,
        64'h00001517_06442483,
        64'h06f42023_16600793,
        64'hdd9ff0ef_51c50513,
        64'h00001517_eadff0ef,
        64'h00090513_00000593,
        64'hdf1ff0ef_52850513,
        64'h00001517_06442903,
        64'h06f42023_10400793,
        64'h20000437_fe079ce3,
        64'hfff78793_00000013,
        64'h04f72023_00a00793,
        64'h20000737_e25ff0ef,
        64'h01212023_00912223,
        64'h00812423_00112623,
        64'h56450513_ff010113,
        64'h00001517_00008067,
        64'h00052503_00008067,
        64'h00b52023_00008067,
        64'h00c68023_fe078ce3,
        64'h0207f793_00074783,
        64'h100006b7_01470713,
        64'h00b68023_10000737,
        64'hfe078ce3_0207f793,
        64'h00074783_100006b7,
        64'h01470713_10000737,
        64'h00074603_0007c583,
        64'h00a787b3_00e78733,
        64'h00455513_e2078793,
        64'h00f57713_00001797,
        64'hfa9ff06f_00f6e7b3,
        64'h00c557b3_00df16b3,
        64'h40ce86b3_00008067,
        64'hfbc61ae3_ff860613,
        64'h00d88023_fe078ce3,
        64'h0207f793_00074783,
        64'h00688023_fe078ce3,
        64'h0207f793_00074783,
        64'h0007c683_0006c303,
        64'h00f807b3_00d806b3,
        64'h00f7f793_0046d693,
        64'h0ff7f693_00f5d7b3,
        64'h0407c863_fe060793,
        64'hff800e13_100008b7,
        64'h01f00e93_03800613,
        64'h01470713_eac80813,
        64'h00159f13_10000737,
        64'h00001817_00008067,
        64'hfa661ee3_ff860613,
        64'h00d80023_fe078ce3,
        64'h0207f793_00074783,
        64'h01180023_fe078ce3,
        64'h0207f793_00074783,
        64'h0007c683_0006c883,
        64'h00f587b3_00d586b3,
        64'h00f7f793_0046d693,
        64'h0ff7f693_00c557b3,
        64'hff800313_10000837,
        64'h01800613_01470713,
        64'hf1458593_10000737,
        64'h00001597_00008067,
        64'h00f58023_0007c783,
        64'h00e580a3_00a787b3,
        64'h00455513_00074703,
        64'h00e78733_f4078793,
        64'h00f57713_00001797,
        64'h00008067_fe0694e3,
        64'h00150513_00154683,
        64'h00d60023_fe078ce3,
        64'h0207f793_00074783,
        64'h10000637_01470713,
        64'h10000737_02068663,
        64'h00054683_00008067,
        64'h00b70823_01070423,
        64'h01170623_00a70223,
        64'h0ff57513_01c70023,
        64'h00855513_0ff57e13,
        64'h02000593_fc700813,
        64'h00300893_00d70623,
        64'hf8000693_00070223,
        64'h10000737_02b55533,
        64'h00459593_00008067,
        64'h00a68023_fe078ce3,
        64'h0207f793_00074783,
        64'h100006b7_01470713,
        64'h10000737_00008067,
        64'h02057513_0147c503,
        64'h100007b7_00008067,
        64'h00054503_00008067,
        64'h00b50023_00008067,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_800004b7,
        64'h18858593_00001597,
        64'hf1402573_ff24c6e3,
        64'h40090913_02000937,
        64'h00448493_fe091ee3,
        64'h0004a903_00092023,
        64'h00990933_00291913,
        64'hf1402973_020004b7,
        64'hfe090ae3_00897913,
        64'h34402973_10500073,
        64'hff24c6e3_40090913,
        64'h02000937_00448493,
        64'h0124a023_00100913,
        64'h020004b7_038010ef,
        64'h84000137_03249463,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
